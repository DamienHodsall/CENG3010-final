library ieee;
use ieee.std_logic_1164;
use ieee.numeric_bit;

entity password is
    port (
        keypress : in std_logic;
        key : in std_logic_vector(0 to 3);
        
         )
